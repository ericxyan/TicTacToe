module TicTacToe(
//	Clock Input
  input CLOCK_50,	//	50 MHz
  input CLOCK_27,     //      27 MHz
//	Push Button
  input [3:0] KEY,      //	Pushbutton[3:0]
//	DPDT Switch
  input [17:0] SW,		//	Toggle Switch[17:0]
//	7-SEG Display
  output [6:0]	HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7,  // Seven Segment Digits
//	LED
  output [8:0]	LEDG,  //	LED Green[8:0]
  output [17:0] LEDR,  //	LED Red[17:0]
//	GPIO
 inout [35:0] GPIO_0,GPIO_1,	//	GPIO Connections
//	TV Decoder
//TD_DATA,    	//	TV Decoder Data bus 8 bits
//TD_HS,		//	TV Decoder H_SYNC
//TD_VS,		//	TV Decoder V_SYNC
  output TD_RESET,	//	TV Decoder Reset
// VGA
  output VGA_CLK,   						//	VGA Clock
  output VGA_HS,							//	VGA H_SYNC
  output VGA_VS,							//	VGA V_SYNC
  output VGA_BLANK,						//	VGA BLANK
  output VGA_SYNC,						//	VGA SYNC
  output [9:0] VGA_R,   						//	VGA Red[9:0]
  output [9:0] VGA_G,	 						//	VGA Green[9:0]
  output [9:0] VGA_B   						//	VGA Blue[9:0]
);

//	All inout port turn to tri-state
assign	GPIO_0		=	36'hzzzzzzzzz;
assign	GPIO_1		=	36'hzzzzzzzzz;

wire RST;
assign RST = KEY[0];

// reset delay gives some time for peripherals to initialize
wire DLY_RST;
Reset_Delay r0(	.iCLK(CLOCK_50),.oRESET(DLY_RST) );

// Send switches to red leds 
assign LEDR = SW;

// Turn off green leds
assign LEDG = 8'h00;

wire [6:0] blank = 7'b111_1111;

// blank unused 7-segment digits
assign HEX0 = blank;
assign HEX1 = blank;
assign HEX2 = blank;
assign HEX3 = blank;
assign HEX4 = blank;
assign HEX5 = blank;
assign HEX6 = blank;
assign HEX7 = blank;

wire		VGA_CTRL_CLK;
wire		AUD_CTRL_CLK;
wire [9:0]	mVGA_R;
wire [9:0]	mVGA_G;
wire [9:0]	mVGA_B;
wire [9:0]	mCoord_X;
wire [9:0]	mCoord_Y;

assign	TD_RESET = 1'b1; // Enable 27 MHz

VGA_Audio_PLL 	p1 (	
	.areset(~DLY_RST),
	.inclk0(CLOCK_27),
	.c0(VGA_CTRL_CLK),
	.c1(AUD_CTRL_CLK),
	.c2(VGA_CLK)
);


// Cursor
reg [9:0] cursor_x = 70;
reg [9:0] cursor_y = 70;

/* Square
	sqaure[21:12]: x
	square[11:2]: y
	square[1:0]: player
	*/
reg [8:0] square;
reg player = 1;
/**
	SW[0]: Move right. 
	SW[1]: Move left. 
	SW[2]: Move down. 
	SW[3]: Move up. 
*/
always @ (posedge KEY[1]) begin
	// move right
	if(cursor_x < 390 && SW[0])
		cursor_x = cursor_x + 160;
	// move left
	if(cursor_x > 70 && SW[1])
		cursor_x = cursor_x - 160;
	// move down
	if((cursor_y < 390) && SW[2])
		cursor_y = cursor_y + 160;
	// move up
	if((cursor_y > 70) && SW[3])
		cursor_y = cursor_y - 160;
	// Draw
	if(SW[4]) begin
		if(cursor_x == 70 && cursor_y == 70) 
			square[0] = player;
		if(cursor_x == 230 && cursor_y == 70) 
			square[1] = player;
		if(cursor_x == 390 && cursor_y == 70) 
			square[2] = player;
		if(cursor_x == 70 && cursor_y == 230) 
			square[3] = player;
		if(cursor_x == 230 && cursor_y == 230) 
			square[4] = player;
		if(cursor_x == 390 && cursor_y ==230) 
			square[5] = player;
		if(cursor_x == 70 && cursor_y == 390) 
			square[6] = player;
		if(cursor_x == 230 && cursor_y == 390) 
			square[7] = player;
		if(cursor_x == 390 && cursor_y == 390) 
			square[8] = player;
		if(player == 1)
			player = 2;
		else
			player = 1;
	end
end


wire [9:0] r, g, b;

// Board
board c1(mCoord_X, mCoord_Y, cursor_x, cursor_y, square, r, g, b);

assign mVGA_R = r;
assign mVGA_G = g;
assign mVGA_B = b;

/*
VGA_Controller	u1 (	
// Host Side
	.iCursor_RGB_EN(4'h7),
	.iRed(mVGA_R),
	.iGreen(mVGA_G),
	.iBlue(mVGA_B),
	.oCoord_X(mCoord_X),
	.oCoord_Y(mCoord_Y),
//  VGA Side
	.oVGA_R(VGA_R),
	.oVGA_G(VGA_G),
	.oVGA_B(VGA_B),
	.oVGA_H_SYNC(VGA_HS),
	.oVGA_V_SYNC(VGA_VS),
	.oVGA_SYNC(VGA_SYNC),
	.oVGA_BLANK(VGA_BLANK),
//   Control Signal
	.iCLK(VGA_CTRL_CLK),
	.iRST_N(DLY_RST&KEY[0])	
);
*/


vga_sync u1(
   .iCLK(VGA_CTRL_CLK),
   .iRST_N(DLY_RST&KEY[0]),	
   .iRed(mVGA_R),
   .iGreen(mVGA_G),
   .iBlue(mVGA_B),
   // pixel coordinates
   .px(mCoord_X),
   .py(mCoord_Y),
   // VGA Side
   .VGA_R(VGA_R),
   .VGA_G(VGA_G),
   .VGA_B(VGA_B),
   .VGA_H_SYNC(VGA_HS),
   .VGA_V_SYNC(VGA_VS),
   .VGA_SYNC(VGA_SYNC),
   .VGA_BLANK(VGA_BLANK)
);


endmodule